				when "00000000000000000000000000000000" => START_BRAM_dout <= "11111111111111111111111111111110";
				when "00000000000000000000000000000100" => START_BRAM_dout <= "00000000000000000000000000000000";
				when "00000000000000000000000000001000" => START_BRAM_dout <= "00000000000000000000000000000010";
				when "00000000000000000000000000001100" => START_BRAM_dout <= "00000000000000000000000000000101";
				when "00000000000000000000000000010000" => START_BRAM_dout <= "00000000000000000000000000000101";
				when "00000000000000000000000000010100" => START_BRAM_dout <= "00000000000000000000000000001000";
				when "00000000000000000000000000011000" => START_BRAM_dout <= "00000000000000000000000000001000";
				when "00000000000000000000000000011100" => START_BRAM_dout <= "00000000000000000000000000001011";
				when "00000000000000000000000000100000" => START_BRAM_dout <= "00000000000000000000000000001011";
				when "00000000000000000000000000100100" => START_BRAM_dout <= "00000000000000000000000000001110";
				when "00000000000000000000000000101000" => START_BRAM_dout <= "00000000000000000000000000001111";
				when "00000000000000000000000000101100" => START_BRAM_dout <= "00000000000000000000000000010010";
				when "00000000000000000000000000110000" => START_BRAM_dout <= "00000000000000000000000000001111";
				when "00000000000000000000000000110100" => START_BRAM_dout <= "00000000000000000000000000001111";
				when "00000000000000000000000000111000" => START_BRAM_dout <= "00000000000000000000000000010010";
				when "00000000000000000000000000111100" => START_BRAM_dout <= "00000000000000000000000000010010";
				when "00000000000000000000000001000000" => START_BRAM_dout <= "00000000000000000000000000010101";
				when "00000000000000000000000001000100" => START_BRAM_dout <= "00000000000000000000000000010110";
				when "00000000000000000000000001001000" => START_BRAM_dout <= "00000000000000000000000000010111";
				when "00000000000000000000000001001100" => START_BRAM_dout <= "00000000000000000000000000011000";
				when "00000000000000000000000001010000" => START_BRAM_dout <= "00000000000000000000000000011001";
				when "00000000000000000000000001010100" => START_BRAM_dout <= "00000000000000000000000000011001";
				when "00000000000000000000000001011000" => START_BRAM_dout <= "00000000000000000000000000011100";
				when "00000000000000000000000001011100" => START_BRAM_dout <= "00000000000000000000000000011100";
