				when "00000000000000000000000000000000" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000000000100" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000000001000" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000000001100" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000000010000" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000000010100" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000000011000" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000000011100" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000000100000" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000000100100" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000000101000" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000000101100" => NB_BRAM_dout <= "00000000000000000000000000000001";
				when "00000000000000000000000000110000" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000000110100" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000000111000" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000000111100" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000001000000" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000001000100" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000001001000" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000001001100" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000001010000" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000001010100" => NB_BRAM_dout <= "00000000000000000000000011100000";
				when "00000000000000000000000001011000" => NB_BRAM_dout <= "00000000000000000000000100100000";
				when "00000000000000000000000001011100" => NB_BRAM_dout <= "00000000000000000000000011100000";
