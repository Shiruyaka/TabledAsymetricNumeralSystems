				when "00000000000000000000000000000000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000110111";
				when "00000000000000000000000000000100" => ENCODING_TABLE_BRAM_dout <= "00110010001100100011001000110011";
				when "00000000000000000000000000001000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000100101";
				when "00000000000000000000000000001100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000101110";
				when "00000000000000000000000000010000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000110011";
				when "00000000000000000000000000010100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000111100";
				when "00000000000000000000000000011000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000101010";
				when "00000000000000000000000000011100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000100001";
				when "00000000000000000000000000100000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000111000";
				when "00000000000000000000000000100100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000101111";
				when "00000000000000000000000000101000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000100110";
				when "00000000000000000000000000101100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000111101";
				when "00000000000000000000000000110000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000110100";
				when "00000000000000000000000000110100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000100010";
				when "00000000000000000000000000111000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000101011";
				when "00000000000000000000000000111100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000111001";
				when "00000000000000000000000001000000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000110000";
				when "00000000000000000000000001000100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000110101";
				when "00000000000000000000000001001000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000111110";
				when "00000000000000000000000001001100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000101100";
				when "00000000000000000000000001010000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000100011";
				when "00000000000000000000000001010100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000111010";
				when "00000000000000000000000001011000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000110001";
				when "00000000000000000000000001011100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000101000";
				when "00000000000000000000000001100000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000111111";
				when "00000000000000000000000001100100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000110110";
				when "00000000000000000000000001101000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000101101";
				when "00000000000000000000000001101100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000100100";
				when "00000000000000000000000001110000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000111011";
				when "00000000000000000000000001110100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000110010";
				when "00000000000000000000000001111000" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000100000";
				when "00000000000000000000000001111100" => ENCODING_TABLE_BRAM_dout <= "00000000000000000000000000101001";
